module mem(
	
	input clk,
	
	output SCL,
	inout SDA
	
	
);



endmodule


